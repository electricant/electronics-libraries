.MODEL 10bq040 d
+IS=2.13126e-05 RS=0.123203 N=1.53952 EG=0.600841
+XTI=3.78803 BV=40 IBV=0.0001 CJO=1.53747e-10
+VJ=1.5 M=0.476132 FC=0.5 TT=0
+KF=0 AF=1
* Model generated on May 28, 96
* Model format: SPICE3

