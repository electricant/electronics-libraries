.MODEL 20ETS12 d
+IS=8.28224e-09 RS=0.00791517 N=1.61051 EG=1.12793
+XTI=0.5 BV=1000 IBV=0.0001 CJO=1e-11
+VJ=0.7 M=0.5 FC=0.5 TT=1e-09
+KF=0 AF=1
* Model generated on Jan 30, 96
* Model format: SPICE3

